library verilog;
use verilog.vl_types.all;
entity array_multiplier_tb is
end array_multiplier_tb;
