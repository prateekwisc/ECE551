library verilog;
use verilog.vl_types.all;
entity t_MACchange is
end t_MACchange;
