library verilog;
use verilog.vl_types.all;
entity t_MAC is
end t_MAC;
