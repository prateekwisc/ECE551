library verilog;
use verilog.vl_types.all;
entity t_FAGP_1bit is
end t_FAGP_1bit;
