library verilog;
use verilog.vl_types.all;
entity t_PIIR is
end t_PIIR;
