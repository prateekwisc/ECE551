library verilog;
use verilog.vl_types.all;
entity test_booth is
end test_booth;
