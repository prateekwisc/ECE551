library verilog;
use verilog.vl_types.all;
entity t_add3_operator is
end t_add3_operator;
