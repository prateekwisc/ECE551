library verilog;
use verilog.vl_types.all;
entity t_CLA_16bit is
end t_CLA_16bit;
