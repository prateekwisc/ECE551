library verilog;
use verilog.vl_types.all;
entity t_CLU_4bit is
end t_CLU_4bit;
