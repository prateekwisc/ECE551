library verilog;
use verilog.vl_types.all;
entity t_ssp is
end t_ssp;
