library verilog;
use verilog.vl_types.all;
entity t_add3_struct is
end t_add3_struct;
