library verilog;
use verilog.vl_types.all;
entity t_receive is
end t_receive;
