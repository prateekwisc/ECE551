library verilog;
use verilog.vl_types.all;
entity t_booth is
end t_booth;
