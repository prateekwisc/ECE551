library verilog;
use verilog.vl_types.all;
entity t_carry_skip is
end t_carry_skip;
