library verilog;
use verilog.vl_types.all;
entity t_errors is
end t_errors;
