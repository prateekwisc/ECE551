library verilog;
use verilog.vl_types.all;
entity t_transmit is
end t_transmit;
